module Adder(input [31:0] A, B, output reg [31:0] sum);

  assign sum = A + B;

endmodule
