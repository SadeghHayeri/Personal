<<<<<<< HEAD
module Adder(input [31:0] A, B, output [31:0] sum);
=======
module Adder(input [31:0] A, B, output reg [31:0] sum);

>>>>>>> 2d3cf3cc6908a26a8f298864c55aedea620bf858
  assign sum = A + B;
endmodule
